library IEEE;
use IEEE.STD_LOGIC_1164.all;


package Basys2 is

	subtype LcdDigit is std_logic_vector(7 downto 0);	
	type LcdDigits is array(3 downto 0) of LcdDigit;	

end Basys2;

package body Basys2 is
end Basys2;

